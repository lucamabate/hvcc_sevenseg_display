magic
tech sky130A
magscale 1 2
timestamp 1669817923
<< obsli1 >>
rect 236104 340159 413848 455521
<< obsm1 >>
rect 2958 6808 580782 703044
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 2962 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580778 703610
rect 2962 6423 580778 703464
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 697140 583440 697237
rect 246 697004 583440 697140
rect 246 684484 583586 697004
rect 560 684084 583586 684484
rect 246 684076 583586 684084
rect 246 683676 583440 684076
rect 246 671428 583586 683676
rect 560 671028 583586 671428
rect 246 670884 583586 671028
rect 246 670484 583440 670884
rect 246 658372 583586 670484
rect 560 657972 583586 658372
rect 246 657556 583586 657972
rect 246 657156 583440 657556
rect 246 645316 583586 657156
rect 560 644916 583586 645316
rect 246 644228 583586 644916
rect 246 643828 583440 644228
rect 246 632260 583586 643828
rect 560 631860 583586 632260
rect 246 631036 583586 631860
rect 246 630636 583440 631036
rect 246 619340 583586 630636
rect 560 618940 583586 619340
rect 246 617708 583586 618940
rect 246 617308 583440 617708
rect 246 606284 583586 617308
rect 560 605884 583586 606284
rect 246 604380 583586 605884
rect 246 603980 583440 604380
rect 246 593228 583586 603980
rect 560 592828 583586 593228
rect 246 591188 583586 592828
rect 246 590788 583440 591188
rect 246 580172 583586 590788
rect 560 579772 583586 580172
rect 246 577860 583586 579772
rect 246 577460 583440 577860
rect 246 567116 583586 577460
rect 560 566716 583586 567116
rect 246 564532 583586 566716
rect 246 564132 583440 564532
rect 246 554060 583586 564132
rect 560 553660 583586 554060
rect 246 551340 583586 553660
rect 246 550940 583440 551340
rect 246 541004 583586 550940
rect 560 540604 583586 541004
rect 246 538012 583586 540604
rect 246 537612 583440 538012
rect 246 528084 583586 537612
rect 560 527684 583586 528084
rect 246 524684 583586 527684
rect 246 524284 583440 524684
rect 246 515028 583586 524284
rect 560 514628 583586 515028
rect 246 511492 583586 514628
rect 246 511092 583440 511492
rect 246 501972 583586 511092
rect 560 501572 583586 501972
rect 246 498164 583586 501572
rect 246 497764 583440 498164
rect 246 488916 583586 497764
rect 560 488516 583586 488916
rect 246 484836 583586 488516
rect 246 484436 583440 484836
rect 246 475860 583586 484436
rect 560 475460 583586 475860
rect 246 471644 583586 475460
rect 246 471244 583440 471644
rect 246 462804 583586 471244
rect 560 462404 583586 462804
rect 246 458316 583586 462404
rect 246 457916 583440 458316
rect 246 449748 583586 457916
rect 560 449348 583586 449748
rect 246 444988 583586 449348
rect 246 444588 583440 444988
rect 246 436828 583586 444588
rect 560 436428 583586 436828
rect 246 431796 583586 436428
rect 246 431396 583440 431796
rect 246 423772 583586 431396
rect 560 423372 583586 423772
rect 246 418468 583586 423372
rect 246 418068 583440 418468
rect 246 410716 583586 418068
rect 560 410316 583586 410716
rect 246 405140 583586 410316
rect 246 404740 583440 405140
rect 246 397660 583586 404740
rect 560 397260 583586 397660
rect 246 391948 583586 397260
rect 246 391548 583440 391948
rect 246 384604 583586 391548
rect 560 384204 583586 384604
rect 246 378620 583586 384204
rect 246 378220 583440 378620
rect 246 371548 583586 378220
rect 560 371148 583586 371548
rect 246 365292 583586 371148
rect 246 364892 583440 365292
rect 246 358628 583586 364892
rect 560 358228 583586 358628
rect 246 352100 583586 358228
rect 246 351700 583440 352100
rect 246 345572 583586 351700
rect 560 345172 583586 345572
rect 246 338772 583586 345172
rect 246 338372 583440 338772
rect 246 332516 583586 338372
rect 560 332116 583586 332516
rect 246 325444 583586 332116
rect 246 325044 583440 325444
rect 246 319460 583586 325044
rect 560 319060 583586 319460
rect 246 312252 583586 319060
rect 246 311852 583440 312252
rect 246 306404 583586 311852
rect 560 306004 583586 306404
rect 246 298924 583586 306004
rect 246 298524 583440 298924
rect 246 293348 583586 298524
rect 560 292948 583586 293348
rect 246 285596 583586 292948
rect 246 285196 583440 285596
rect 246 280292 583586 285196
rect 560 279892 583586 280292
rect 246 272404 583586 279892
rect 246 272004 583440 272404
rect 246 267372 583586 272004
rect 560 266972 583586 267372
rect 246 259076 583586 266972
rect 246 258676 583440 259076
rect 246 254316 583586 258676
rect 560 253916 583586 254316
rect 246 245748 583586 253916
rect 246 245348 583440 245748
rect 246 241260 583586 245348
rect 560 240860 583586 241260
rect 246 232556 583586 240860
rect 246 232156 583440 232556
rect 246 228204 583586 232156
rect 560 227804 583586 228204
rect 246 219228 583586 227804
rect 246 218828 583440 219228
rect 246 215148 583586 218828
rect 560 214748 583586 215148
rect 246 205900 583586 214748
rect 246 205500 583440 205900
rect 246 202092 583586 205500
rect 560 201692 583586 202092
rect 246 192708 583586 201692
rect 246 192308 583440 192708
rect 246 189036 583586 192308
rect 560 188636 583586 189036
rect 246 179380 583586 188636
rect 246 178980 583440 179380
rect 246 176116 583586 178980
rect 560 175716 583586 176116
rect 246 166052 583586 175716
rect 246 165652 583440 166052
rect 246 163060 583586 165652
rect 560 162660 583586 163060
rect 246 152860 583586 162660
rect 246 152460 583440 152860
rect 246 150004 583586 152460
rect 560 149604 583586 150004
rect 246 139532 583586 149604
rect 246 139132 583440 139532
rect 246 136948 583586 139132
rect 560 136548 583586 136948
rect 246 126204 583586 136548
rect 246 125804 583440 126204
rect 246 113012 583586 125804
rect 246 112612 583440 113012
rect 246 110836 583586 112612
rect 560 110436 583586 110836
rect 246 99684 583586 110436
rect 246 99284 583440 99684
rect 246 97780 583586 99284
rect 560 97380 583586 97780
rect 246 86356 583586 97380
rect 246 85956 583440 86356
rect 246 84860 583586 85956
rect 560 84460 583586 84860
rect 246 73164 583586 84460
rect 246 72764 583440 73164
rect 246 71804 583586 72764
rect 560 71404 583586 71804
rect 246 59836 583586 71404
rect 246 59436 583440 59836
rect 246 58748 583586 59436
rect 560 58348 583586 58748
rect 246 46508 583586 58348
rect 246 46108 583440 46508
rect 246 45692 583586 46108
rect 560 45292 583586 45692
rect 246 33316 583586 45292
rect 246 32916 583440 33316
rect 246 32636 583586 32916
rect 560 32236 583586 32636
rect 246 19988 583586 32236
rect 246 19588 583440 19988
rect 246 19580 583586 19588
rect 560 19180 583586 19580
rect 246 6796 583586 19180
rect 246 6660 583440 6796
rect 560 6427 583440 6660
<< metal4 >>
rect -23776 -22704 -23156 726640
rect -20666 -19594 -20046 723530
rect -17556 -16484 -16936 720420
rect -14446 -13374 -13826 717310
rect -11336 -10264 -10716 714200
rect -8226 -7154 -7606 711090
rect -5116 -4044 -4496 707980
rect -2006 -934 -1386 704870
rect 1794 -22704 2414 726640
rect 5514 -22704 6134 726640
rect 9234 -22704 9854 726640
rect 12954 -22704 13574 726640
rect 16674 -22704 17294 726640
rect 20394 -22704 21014 726640
rect 24114 -22704 24734 726640
rect 27834 -22704 28454 726640
rect 37794 -22704 38414 726640
rect 41514 -22704 42134 726640
rect 45234 -22704 45854 726640
rect 48954 -22704 49574 726640
rect 52674 -22704 53294 726640
rect 56394 -22704 57014 726640
rect 60114 -22704 60734 726640
rect 63834 -22704 64454 726640
rect 73794 -22704 74414 726640
rect 77514 -22704 78134 726640
rect 81234 -22704 81854 726640
rect 84954 -22704 85574 726640
rect 88674 -22704 89294 726640
rect 92394 -22704 93014 726640
rect 96114 -22704 96734 726640
rect 99834 -22704 100454 726640
rect 109794 -22704 110414 726640
rect 113514 -22704 114134 726640
rect 117234 -22704 117854 726640
rect 120954 -22704 121574 726640
rect 124674 -22704 125294 726640
rect 128394 -22704 129014 726640
rect 132114 -22704 132734 726640
rect 135834 -22704 136454 726640
rect 145794 -22704 146414 726640
rect 149514 -22704 150134 726640
rect 153234 -22704 153854 726640
rect 156954 -22704 157574 726640
rect 160674 -22704 161294 726640
rect 164394 -22704 165014 726640
rect 168114 -22704 168734 726640
rect 171834 -22704 172454 726640
rect 181794 -22704 182414 726640
rect 185514 -22704 186134 726640
rect 189234 -22704 189854 726640
rect 192954 -22704 193574 726640
rect 196674 -22704 197294 726640
rect 200394 -22704 201014 726640
rect 204114 -22704 204734 726640
rect 207834 -22704 208454 726640
rect 217794 -22704 218414 726640
rect 221514 -22704 222134 726640
rect 225234 -22704 225854 726640
rect 228954 -22704 229574 726640
rect 232674 -22704 233294 726640
rect 236394 -22704 237014 726640
rect 240114 -22704 240734 726640
rect 243834 -22704 244454 726640
rect 253794 -22704 254414 726640
rect 257514 -22704 258134 726640
rect 261234 -22704 261854 726640
rect 264954 -22704 265574 726640
rect 268674 -22704 269294 726640
rect 272394 -22704 273014 726640
rect 276114 -22704 276734 726640
rect 279834 -22704 280454 726640
rect 289794 -22704 290414 726640
rect 293514 -22704 294134 726640
rect 297234 -22704 297854 726640
rect 300954 457612 301574 726640
rect 300954 -22704 301574 338068
rect 304674 -22704 305294 726640
rect 308394 -22704 309014 726640
rect 312114 -22704 312734 726640
rect 315834 457612 316454 726640
rect 315834 -22704 316454 338068
rect 325794 -22704 326414 726640
rect 329514 -22704 330134 726640
rect 333234 -22704 333854 726640
rect 336954 -22704 337574 726640
rect 340674 -22704 341294 726640
rect 344394 -22704 345014 726640
rect 348114 -22704 348734 726640
rect 351834 -22704 352454 726640
rect 361794 457612 362414 726640
rect 361794 -22704 362414 338068
rect 365514 -22704 366134 726640
rect 369234 -22704 369854 726640
rect 372954 -22704 373574 726640
rect 376674 -22704 377294 726640
rect 380394 -22704 381014 726640
rect 384114 -22704 384734 726640
rect 387834 -22704 388454 726640
rect 397794 -22704 398414 726640
rect 401514 -22704 402134 726640
rect 405234 -22704 405854 726640
rect 408954 -22704 409574 726640
rect 412674 -22704 413294 726640
rect 416394 -22704 417014 726640
rect 420114 -22704 420734 726640
rect 423834 -22704 424454 726640
rect 433794 -22704 434414 726640
rect 437514 -22704 438134 726640
rect 441234 -22704 441854 726640
rect 444954 -22704 445574 726640
rect 448674 -22704 449294 726640
rect 452394 -22704 453014 726640
rect 456114 -22704 456734 726640
rect 459834 -22704 460454 726640
rect 469794 -22704 470414 726640
rect 473514 -22704 474134 726640
rect 477234 -22704 477854 726640
rect 480954 -22704 481574 726640
rect 484674 -22704 485294 726640
rect 488394 -22704 489014 726640
rect 492114 -22704 492734 726640
rect 495834 -22704 496454 726640
rect 505794 -22704 506414 726640
rect 509514 -22704 510134 726640
rect 513234 -22704 513854 726640
rect 516954 -22704 517574 726640
rect 520674 -22704 521294 726640
rect 524394 -22704 525014 726640
rect 528114 -22704 528734 726640
rect 531834 -22704 532454 726640
rect 541794 -22704 542414 726640
rect 545514 -22704 546134 726640
rect 549234 -22704 549854 726640
rect 552954 -22704 553574 726640
rect 556674 -22704 557294 726640
rect 560394 -22704 561014 726640
rect 564114 -22704 564734 726640
rect 567834 -22704 568454 726640
rect 577794 -22704 578414 726640
rect 581514 -22704 582134 726640
rect 585310 -934 585930 704870
rect 588420 -4044 589040 707980
rect 591530 -7154 592150 711090
rect 594640 -10264 595260 714200
rect 597750 -13374 598370 717310
rect 600860 -16484 601480 720420
rect 603970 -19594 604590 723530
rect 607080 -22704 607700 726640
<< obsm4 >>
rect 239208 57971 240034 460325
rect 240814 57971 243754 460325
rect 244534 57971 253714 460325
rect 254494 57971 257434 460325
rect 258214 57971 261154 460325
rect 261934 57971 264874 460325
rect 265654 57971 268594 460325
rect 269374 57971 272314 460325
rect 273094 57971 276034 460325
rect 276814 57971 279754 460325
rect 280534 57971 289714 460325
rect 290494 57971 293434 460325
rect 294214 57971 297154 460325
rect 297934 457532 300874 460325
rect 301654 457532 304594 460325
rect 297934 338148 304594 457532
rect 297934 57971 300874 338148
rect 301654 57971 304594 338148
rect 305374 57971 308314 460325
rect 309094 57971 312034 460325
rect 312814 457532 315754 460325
rect 316534 457532 325714 460325
rect 312814 338148 325714 457532
rect 312814 57971 315754 338148
rect 316534 57971 325714 338148
rect 326494 57971 329434 460325
rect 330214 57971 333154 460325
rect 333934 57971 336874 460325
rect 337654 57971 340594 460325
rect 341374 57971 344314 460325
rect 345094 57971 348034 460325
rect 348814 57971 351754 460325
rect 352534 457532 361714 460325
rect 362494 457532 365434 460325
rect 352534 338148 365434 457532
rect 352534 57971 361714 338148
rect 362494 57971 365434 338148
rect 366214 57971 369154 460325
rect 369934 57971 372874 460325
rect 373654 57971 376594 460325
rect 377374 57971 380314 460325
rect 381094 57971 384034 460325
rect 384814 57971 387754 460325
rect 388534 57971 397714 460325
rect 398494 57971 401434 460325
rect 402214 57971 405154 460325
rect 405934 57971 408874 460325
rect 409654 57971 411365 460325
<< metal5 >>
rect -23776 726020 607700 726640
rect -20666 722910 604590 723530
rect -17556 719800 601480 720420
rect -14446 716690 598370 717310
rect -11336 713580 595260 714200
rect -8226 710470 592150 711090
rect -5116 707360 589040 707980
rect -2006 704250 585930 704870
rect -23776 698026 607700 698646
rect -23776 694306 607700 694926
rect -23776 690586 607700 691206
rect -23776 686866 607700 687486
rect -23776 676906 607700 677526
rect -23776 673186 607700 673806
rect -23776 669466 607700 670086
rect -23776 665746 607700 666366
rect -23776 662026 607700 662646
rect -23776 658306 607700 658926
rect -23776 654586 607700 655206
rect -23776 650866 607700 651486
rect -23776 640906 607700 641526
rect -23776 637186 607700 637806
rect -23776 633466 607700 634086
rect -23776 629746 607700 630366
rect -23776 626026 607700 626646
rect -23776 622306 607700 622926
rect -23776 618586 607700 619206
rect -23776 614866 607700 615486
rect -23776 604906 607700 605526
rect -23776 601186 607700 601806
rect -23776 597466 607700 598086
rect -23776 593746 607700 594366
rect -23776 590026 607700 590646
rect -23776 586306 607700 586926
rect -23776 582586 607700 583206
rect -23776 578866 607700 579486
rect -23776 568906 607700 569526
rect -23776 565186 607700 565806
rect -23776 561466 607700 562086
rect -23776 557746 607700 558366
rect -23776 554026 607700 554646
rect -23776 550306 607700 550926
rect -23776 546586 607700 547206
rect -23776 542866 607700 543486
rect -23776 532906 607700 533526
rect -23776 529186 607700 529806
rect -23776 525466 607700 526086
rect -23776 521746 607700 522366
rect -23776 518026 607700 518646
rect -23776 514306 607700 514926
rect -23776 510586 607700 511206
rect -23776 506866 607700 507486
rect -23776 496906 607700 497526
rect -23776 493186 607700 493806
rect -23776 489466 607700 490086
rect -23776 485746 607700 486366
rect -23776 482026 607700 482646
rect -23776 478306 607700 478926
rect -23776 474586 607700 475206
rect -23776 470866 607700 471486
rect -23776 460906 607700 461526
rect -23776 457186 607700 457806
rect -23776 453466 607700 454086
rect -23776 449746 607700 450366
rect -23776 446026 607700 446646
rect -23776 442306 607700 442926
rect -23776 438586 607700 439206
rect -23776 434866 607700 435486
rect -23776 424906 607700 425526
rect -23776 421186 607700 421806
rect -23776 417466 607700 418086
rect -23776 413746 607700 414366
rect -23776 410026 607700 410646
rect -23776 406306 607700 406926
rect -23776 402586 607700 403206
rect -23776 398866 607700 399486
rect -23776 388906 607700 389526
rect -23776 385186 607700 385806
rect -23776 381466 607700 382086
rect -23776 377746 607700 378366
rect -23776 374026 607700 374646
rect -23776 370306 607700 370926
rect -23776 366586 607700 367206
rect -23776 362866 607700 363486
rect -23776 352906 607700 353526
rect -23776 349186 607700 349806
rect -23776 345466 607700 346086
rect -23776 341746 607700 342366
rect -23776 338026 607700 338646
rect -23776 334306 607700 334926
rect -23776 330586 607700 331206
rect -23776 326866 607700 327486
rect -23776 316906 607700 317526
rect -23776 313186 607700 313806
rect -23776 309466 607700 310086
rect -23776 305746 607700 306366
rect -23776 302026 607700 302646
rect -23776 298306 607700 298926
rect -23776 294586 607700 295206
rect -23776 290866 607700 291486
rect -23776 280906 607700 281526
rect -23776 277186 607700 277806
rect -23776 273466 607700 274086
rect -23776 269746 607700 270366
rect -23776 266026 607700 266646
rect -23776 262306 607700 262926
rect -23776 258586 607700 259206
rect -23776 254866 607700 255486
rect -23776 244906 607700 245526
rect -23776 241186 607700 241806
rect -23776 237466 607700 238086
rect -23776 233746 607700 234366
rect -23776 230026 607700 230646
rect -23776 226306 607700 226926
rect -23776 222586 607700 223206
rect -23776 218866 607700 219486
rect -23776 208906 607700 209526
rect -23776 205186 607700 205806
rect -23776 201466 607700 202086
rect -23776 197746 607700 198366
rect -23776 194026 607700 194646
rect -23776 190306 607700 190926
rect -23776 186586 607700 187206
rect -23776 182866 607700 183486
rect -23776 172906 607700 173526
rect -23776 169186 607700 169806
rect -23776 165466 607700 166086
rect -23776 161746 607700 162366
rect -23776 158026 607700 158646
rect -23776 154306 607700 154926
rect -23776 150586 607700 151206
rect -23776 146866 607700 147486
rect -23776 136906 607700 137526
rect -23776 133186 607700 133806
rect -23776 129466 607700 130086
rect -23776 125746 607700 126366
rect -23776 122026 607700 122646
rect -23776 118306 607700 118926
rect -23776 114586 607700 115206
rect -23776 110866 607700 111486
rect -23776 100906 607700 101526
rect -23776 97186 607700 97806
rect -23776 93466 607700 94086
rect -23776 89746 607700 90366
rect -23776 86026 607700 86646
rect -23776 82306 607700 82926
rect -23776 78586 607700 79206
rect -23776 74866 607700 75486
rect -23776 64906 607700 65526
rect -23776 61186 607700 61806
rect -23776 57466 607700 58086
rect -23776 53746 607700 54366
rect -23776 50026 607700 50646
rect -23776 46306 607700 46926
rect -23776 42586 607700 43206
rect -23776 38866 607700 39486
rect -23776 28906 607700 29526
rect -23776 25186 607700 25806
rect -23776 21466 607700 22086
rect -23776 17746 607700 18366
rect -23776 14026 607700 14646
rect -23776 10306 607700 10926
rect -23776 6586 607700 7206
rect -23776 2866 607700 3486
rect -2006 -934 585930 -314
rect -5116 -4044 589040 -3424
rect -8226 -7154 592150 -6534
rect -11336 -10264 595260 -9644
rect -14446 -13374 598370 -12754
rect -17556 -16484 601480 -15864
rect -20666 -19594 604590 -18974
rect -23776 -22704 607700 -22084
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 1794 -22704 2414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 37794 -22704 38414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 73794 -22704 74414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 109794 -22704 110414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 145794 -22704 146414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 181794 -22704 182414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 217794 -22704 218414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 253794 -22704 254414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 289794 -22704 290414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 325794 -22704 326414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 -22704 362414 338068 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 361794 457612 362414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 397794 -22704 398414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 433794 -22704 434414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 469794 -22704 470414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 505794 -22704 506414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 541794 -22704 542414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s 577794 -22704 578414 726640 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 2866 607700 3486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 38866 607700 39486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 74866 607700 75486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 110866 607700 111486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 146866 607700 147486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 182866 607700 183486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 218866 607700 219486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 254866 607700 255486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 290866 607700 291486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 326866 607700 327486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 362866 607700 363486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 398866 607700 399486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 434866 607700 435486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 470866 607700 471486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 506866 607700 507486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 542866 607700 543486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 578866 607700 579486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 614866 607700 615486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 650866 607700 651486 6 vccd1
port 531 nsew power bidirectional
rlabel metal5 s -23776 686866 607700 687486 6 vccd1
port 531 nsew power bidirectional
rlabel metal4 s -8226 -7154 -7606 711090 4 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8226 -7154 592150 -6534 8 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -8226 710470 592150 711090 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 591530 -7154 592150 711090 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 9234 -22704 9854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 45234 -22704 45854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 81234 -22704 81854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 117234 -22704 117854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 153234 -22704 153854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 189234 -22704 189854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 225234 -22704 225854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 261234 -22704 261854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 297234 -22704 297854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 333234 -22704 333854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 369234 -22704 369854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 405234 -22704 405854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 441234 -22704 441854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 477234 -22704 477854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 513234 -22704 513854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s 549234 -22704 549854 726640 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 10306 607700 10926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 46306 607700 46926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 82306 607700 82926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 118306 607700 118926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 154306 607700 154926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 190306 607700 190926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 226306 607700 226926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 262306 607700 262926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 298306 607700 298926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 334306 607700 334926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 370306 607700 370926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 406306 607700 406926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 442306 607700 442926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 478306 607700 478926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 514306 607700 514926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 550306 607700 550926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 586306 607700 586926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 622306 607700 622926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 658306 607700 658926 6 vccd2
port 532 nsew power bidirectional
rlabel metal5 s -23776 694306 607700 694926 6 vccd2
port 532 nsew power bidirectional
rlabel metal4 s -14446 -13374 -13826 717310 4 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -14446 -13374 598370 -12754 8 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -14446 716690 598370 717310 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 597750 -13374 598370 717310 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 16674 -22704 17294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 52674 -22704 53294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 88674 -22704 89294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 124674 -22704 125294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 160674 -22704 161294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 196674 -22704 197294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 232674 -22704 233294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 268674 -22704 269294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 304674 -22704 305294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 340674 -22704 341294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 376674 -22704 377294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 412674 -22704 413294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 448674 -22704 449294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 484674 -22704 485294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 520674 -22704 521294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s 556674 -22704 557294 726640 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 17746 607700 18366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 53746 607700 54366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 89746 607700 90366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 125746 607700 126366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 161746 607700 162366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 197746 607700 198366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 233746 607700 234366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 269746 607700 270366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 305746 607700 306366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 341746 607700 342366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 377746 607700 378366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 413746 607700 414366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 449746 607700 450366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 485746 607700 486366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 521746 607700 522366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 557746 607700 558366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 593746 607700 594366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 629746 607700 630366 6 vdda1
port 533 nsew power bidirectional
rlabel metal5 s -23776 665746 607700 666366 6 vdda1
port 533 nsew power bidirectional
rlabel metal4 s -20666 -19594 -20046 723530 4 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -20666 -19594 604590 -18974 8 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -20666 722910 604590 723530 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 603970 -19594 604590 723530 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 24114 -22704 24734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 60114 -22704 60734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 96114 -22704 96734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 132114 -22704 132734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 168114 -22704 168734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 204114 -22704 204734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 240114 -22704 240734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 276114 -22704 276734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 312114 -22704 312734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 348114 -22704 348734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 384114 -22704 384734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 420114 -22704 420734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 456114 -22704 456734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 492114 -22704 492734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 528114 -22704 528734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 564114 -22704 564734 726640 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 25186 607700 25806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 61186 607700 61806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 97186 607700 97806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 133186 607700 133806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 169186 607700 169806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 205186 607700 205806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 241186 607700 241806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 277186 607700 277806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 313186 607700 313806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 349186 607700 349806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 385186 607700 385806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 421186 607700 421806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 457186 607700 457806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 493186 607700 493806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 529186 607700 529806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 565186 607700 565806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 601186 607700 601806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 637186 607700 637806 6 vdda2
port 534 nsew power bidirectional
rlabel metal5 s -23776 673186 607700 673806 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s -17556 -16484 -16936 720420 4 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -17556 -16484 601480 -15864 8 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -17556 719800 601480 720420 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 600860 -16484 601480 720420 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 20394 -22704 21014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 56394 -22704 57014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 92394 -22704 93014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 128394 -22704 129014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 164394 -22704 165014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 200394 -22704 201014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 236394 -22704 237014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 272394 -22704 273014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 308394 -22704 309014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 344394 -22704 345014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 380394 -22704 381014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 416394 -22704 417014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 452394 -22704 453014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 488394 -22704 489014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 524394 -22704 525014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s 560394 -22704 561014 726640 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 21466 607700 22086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 57466 607700 58086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 93466 607700 94086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 129466 607700 130086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 165466 607700 166086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 201466 607700 202086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 237466 607700 238086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 273466 607700 274086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 309466 607700 310086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 345466 607700 346086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 381466 607700 382086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 417466 607700 418086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 453466 607700 454086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 489466 607700 490086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 525466 607700 526086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 561466 607700 562086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 597466 607700 598086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 633466 607700 634086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal5 s -23776 669466 607700 670086 6 vssa1
port 535 nsew ground bidirectional
rlabel metal4 s -23776 -22704 -23156 726640 4 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 -22704 607700 -22084 8 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 726020 607700 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 607080 -22704 607700 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 27834 -22704 28454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 63834 -22704 64454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 99834 -22704 100454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 135834 -22704 136454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 171834 -22704 172454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 207834 -22704 208454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 243834 -22704 244454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 279834 -22704 280454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 315834 -22704 316454 338068 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 315834 457612 316454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 351834 -22704 352454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 387834 -22704 388454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 423834 -22704 424454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 459834 -22704 460454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 495834 -22704 496454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 531834 -22704 532454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 567834 -22704 568454 726640 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 28906 607700 29526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 64906 607700 65526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 100906 607700 101526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 136906 607700 137526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 172906 607700 173526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 208906 607700 209526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 244906 607700 245526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 280906 607700 281526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 316906 607700 317526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 352906 607700 353526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 388906 607700 389526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 424906 607700 425526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 460906 607700 461526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 496906 607700 497526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 532906 607700 533526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 568906 607700 569526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 604906 607700 605526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 640906 607700 641526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal5 s -23776 676906 607700 677526 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s -5116 -4044 -4496 707980 4 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -5116 -4044 589040 -3424 8 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -5116 707360 589040 707980 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 588420 -4044 589040 707980 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 5514 -22704 6134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 41514 -22704 42134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 77514 -22704 78134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 113514 -22704 114134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 149514 -22704 150134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 185514 -22704 186134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 221514 -22704 222134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 257514 -22704 258134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 293514 -22704 294134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 329514 -22704 330134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 365514 -22704 366134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 401514 -22704 402134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 437514 -22704 438134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 473514 -22704 474134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 509514 -22704 510134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 545514 -22704 546134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s 581514 -22704 582134 726640 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 6586 607700 7206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 42586 607700 43206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 78586 607700 79206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 114586 607700 115206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 150586 607700 151206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 186586 607700 187206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 222586 607700 223206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 258586 607700 259206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 294586 607700 295206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 330586 607700 331206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 366586 607700 367206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 402586 607700 403206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 438586 607700 439206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 474586 607700 475206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 510586 607700 511206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 546586 607700 547206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 582586 607700 583206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 618586 607700 619206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 654586 607700 655206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal5 s -23776 690586 607700 691206 6 vssd1
port 537 nsew ground bidirectional
rlabel metal4 s -11336 -10264 -10716 714200 4 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -11336 -10264 595260 -9644 8 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -11336 713580 595260 714200 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 594640 -10264 595260 714200 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 12954 -22704 13574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 48954 -22704 49574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 84954 -22704 85574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 120954 -22704 121574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 156954 -22704 157574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 192954 -22704 193574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 228954 -22704 229574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 264954 -22704 265574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 300954 -22704 301574 338068 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 300954 457612 301574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 336954 -22704 337574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 372954 -22704 373574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 408954 -22704 409574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 444954 -22704 445574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 480954 -22704 481574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 516954 -22704 517574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal4 s 552954 -22704 553574 726640 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 14026 607700 14646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 50026 607700 50646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 86026 607700 86646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 122026 607700 122646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 158026 607700 158646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 194026 607700 194646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 230026 607700 230646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 266026 607700 266646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 302026 607700 302646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 338026 607700 338646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 374026 607700 374646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 410026 607700 410646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 446026 607700 446646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 482026 607700 482646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 518026 607700 518646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 554026 607700 554646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 590026 607700 590646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 626026 607700 626646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 662026 607700 662646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal5 s -23776 698026 607700 698646 6 vssd2
port 538 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6810516
string GDS_FILE /home/designer-01/designs/hvcc_sevenseg_display/openlane/user_project_wrapper/runs/22_11_30_06_17/results/signoff/user_project_wrapper.magic.gds
string GDS_START 5633078
<< end >>

